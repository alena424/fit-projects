BZh91AY&SY��� �߀Py����߰?���P~t���  �RmL���	�&�h�a��F��`LM&L�LM2100	MjOP �     `LM&L�LM2100	i�zh�M)�xM4�H��FCj0�?P%	*�-H��!3���Q��ZM��1�m/?�D$�K��Q�U��#V��=��aF��}�F-iH��<����-�0l��sS~�v�(�d�:�"�(@KC#9$�h���+��'B���YX��nnX��	��9�59��(�:*xQKE�(�e��de�A��%,G��X�DZ��_�{���|��E1�R�^EfK��E(���F��)�`����}�Єʉ$�Hq7��o65=�z�n�j�T�9��!@��DM��wI�i$��hAFU��`^���E*q $��k��_rh-G��W�k]�3�2tYܽ�n5���OF7�Z>�9! ��c��7�4 ~#�+0�'Q�.�r��?�,�����1,�r*v�{����q��nlD�(�L�+#	���pgJ���$J���!(��-QH�%(V���u�QYm�)��vOz��L�+3��rA��Id���:���~�
�!3��T
O:g�)�¥���̏�J�f!�N4���SZ�L�.����5�����b����d�����r���3�mUMk��0�F��a~�ԌǞ����A�l[�Dhji��ҖT�L6i-�YY>ޤwe��H�x� Zl�}�ԯ�a# �	��$����1�X*����C�L���*-���7�h�6���C*����J� RWU�J]#�j�OfAǱG���y��Ѧ@����-'�0@��Pd(5��9-���Ԓ�6r�לW�9`���M��~��Ӳ��#0uX
��<1���	���n��:�@s�7���E�k������s�2ĩ��M!@�L�Jl����#l�7aUV�#ʥXе)�����8Sh��b&�0L�rE8P����